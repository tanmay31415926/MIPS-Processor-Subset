module instruction_memory (
    input wire [31:0] address,         // PC value
    output wire [31:0] instruction     // Fetched instruction
);

    reg [31:0] memory [0:255];         // 256 words = 1 KB instruction memory

    initial begin
        // Instruction encodings
//        memory[0]  = 32'b100011_00000_00001_0000000000000000;  // lw $1, 0($0)
//        memory[1]  = 32'b100011_00000_00010_0000000000000100;  // lw $2, 4($0)
//        memory[2]  = 32'b100011_00000_00011_0000000000001000;  // lw $3, 8($0)
//        memory[3]  = 32'b000000_00000_00000_00100_00000_100000; // add $4, $0, $0
//        memory[4]  = 32'b100011_00000_00101_0000000000001100;  // lw $5, 12($0)
//        memory[5]  = 32'b000000_00100_00001_00100_00000_100000; // add $4, $4, $1
//        memory[6]  = 32'b000000_00100_00010_00100_00000_100000; // add $4, $4, $2
//        memory[7]  = 32'b000000_00011_00101_00011_00000_100010; // sub $3, $3, $5
//        memory[8] = 32'b101011_00000_00100_0000000110010000;  // sw $4, 400($0)
//        memory[9]  = 32'b000100_00011_00000_0000000000000001;  // beq $3, $0, done (PC+4+1*4 = addr 40)
    
//        memory[10]  = 32'b000100_00000_00000_1111111111111010;  // beq $0, $0, loop (offset = -5)
//        memory[11]  = 32'b000100_00000_00000_1111111111111111;  // beq $0, $0, loop (offset = -1) loop at done
////        memory[10]  = 32'b000010_00000000000000000000000101;  // jumping to instruction 5
        // Load n from memory[0]
        memory[0]  = 32'b100011_00000_00010_0000000000000000; // lw $2, 0($0)      ; n
        memory[1]  = 32'b000000_00000_00000_00011_00000_100000; // add $3, $0, $0    ; first = 0
        memory[2]  = 32'b000000_00000_00001_00100_00000_100000; // add $4, $0, $1    ; second = 1 (use $1 as temp)
        memory[3]  = 32'b000000_00000_00000_00110_00000_100000; // add $6, $0, $0    ; counter = 0
        
        // Label: loop
        memory[4]  = 32'b101011_00001_00011_0000000000000010; // sw $3, 2($1)       ; store first
        memory[5]  = 32'b000000_00011_00100_00101_00000_100000; // add $5, $3, $4    ; next = first + second
        memory[6]  = 32'b000000_00100_00000_00011_00000_100000; // add $3, $4, $0    ; first = second
        memory[7]  = 32'b000000_00101_00000_00100_00000_100000; // add $4, $5, $0    ; second = next
        memory[8]  = 32'b000000_00110_00001_00110_00000_100000; // add $6, $6, $1    ; counter += 1
        memory[9]  = 32'b000000_00110_00000_00111_00000_100000; // add $7, $6, $0    ; temp = counter
        memory[10] = 32'b000000_00111_00010_00111_00000_101010; // slt $7, $7, $2    ; if counter < n
         
        memory[11] = 32'b101011_00000_00100_0000000110010000; // sw $4, 400($0)
        memory[12] = 32'b000100_00111_00001_1111111111111000; // be $7, $1, -8   ; branch to loop (PC-relative)
        memory[13]  = 32'b000100_00000_00000_1111111111111111;  // beq $0, $0, loop (offset = -1) loop at done
        
      

// function fib:
// if n == 0: return 0
    // Initialize $2 and $3 from memory (example: mem[100] and mem[104])
//memory[0] = 32'b100011_00000_00010_0000000001100100; // lw $2, 100($0)
//memory[1] = 32'b100011_00000_00011_0000000001101000; // lw $3, 104($0)
//memory[2] = 32'b000011_00000_00000_0000000000000110; // jal 6 (func starts at memory[6])
//memory[3] = 32'b000000_00000_00000_00000_00000_000000; // nop (optional)
//memory[4] = 32'b101011_00000_00100_0000000001101100; // sw $4, 108($0)
//memory[5] = 32'b000000_00000_00000_00000_00000_000000; // end: nop

//// func:
//memory[6] = 32'b000000_00010_00011_00100_00000_100100; // add $4, $2, $3
//memory[7] = 32'b000000_11111_00000_00000_00000_001000; // jr $31

       
        
    end

    assign instruction = memory[address[9:2]]; // Word aligned access (ignore lower 2 bits)

endmodule
